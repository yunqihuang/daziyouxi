module sec_timer()